entity Dec2_4EnDemo is
 port(SW : std_logic_vector(2 downto 0);
 LEDG : std_logic_vector(3 downto 0));
architecture Shell of Dec2_4EnDemo is
begin
 system_core : work entity.Dec2_4En(BehavEquations)
 port map(enable <= SW(2);
 inputs <= SW;
 outputs => LEDG(3 downto 0);
end Dec2_4EnDemo; 