library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity SeqShiftUnit is
	port(clk : in std_logic;   -- clock 
		  dataIn : in std_logic_vector(7 downto 0); -- input com 8 bits
		  siLeft : in std_logic;       -- esquerda
		  siRight : in std_logic;      -- direita 
		  loadEn : in std_logic;
		  rotate : in std_logic;
		  dirLeft : in std_logic;
        shArith : in std_logic;
        dataOut : out std_logic_vector(7 downto 0)); -- output com 8 bits 
end SeqShiftUnit;

architecture Behavioral of SeqShiftUnit is
 signal s_shiftReg : std_logic_vector(7 downto 0);    

 begin
  process(clk)
 begin
 if (falling_edge(clk)) then   -- clock v
 -- paralel load
 if (loadEn = '1') then
 s_shiftReg <= dataIn;
 
 -- rotate 
 elsif (rotate = '1') then
 if (dirLeft = '1') then
 s_shiftReg <= s_shiftReg(6 downto 0) & s_shiftReg(7);
 else
 s_shiftReg <= s_shiftReg(0) & s_shiftReg(7 downto 1);
 end if;
 
 -- shifts aritmeticos
 elsif (shArith = '1') then
   -- shift left
	if ( dirLeft = '1') then 
	 s_shiftReg <= s_shiftReg(6 downto 0) & '0';
	-- shift right
	else
	s_shiftReg <= s_shiftReg(7) & s_shiftReg(7 downto 1);
	end if;
-- shifts logicos 
  else
	--Shift Left
	 if (dirLeft = '1') then
		s_shiftReg <= s_shiftReg(6 downto 0) & siLeft;
	--Shift Right
	 else	
	   s_shiftReg <= siRight & s_shiftReg(7 downto 1);
 end if; 
 end if;
 end if;
 end process;
 dataOut <= s_shiftReg;
end Behavioral; 